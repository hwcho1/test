������� �����͸� pull�ϱ� ���� �Ἥ push�Ϸ��� �ؽ�Ʈ����
