asdjhgslkj
qqq
www
eee
+rrr
@DDD
+ttt
1234
dfsdfsdsdfsfddfsdfsdfsdfsdfsdf
+sfsdfsdf+erer
+werwerwr
