qqq
www
eee
+rrr
@DDD
+ttt
1234
