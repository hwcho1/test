qqq
www
eee
+rrr
