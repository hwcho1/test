int a
class
int b
int c
int d;
