qqq
www
eee
+rrr
@DDD
