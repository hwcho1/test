class
	rand logic [3:0] a;
	rand logic [3:0] b;

endclass
