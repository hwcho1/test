logic a
logic b
