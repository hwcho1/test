qqq
www
eee
+rrr
@DDD
+ttt
